* C:\Users\Pc\Documents\CS_LAB_Spise\lab13.sch

* Schematics Version 9.1 - Web Update 1
* Wed Aug 05 18:46:15 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "lab13.net"
.INC "lab13.als"


.probe


.END
