* C:\Users\Pc\Documents\CS_LAB_Spise\complex_matlab_analysis.sch

* Schematics Version 9.1 - Web Update 1
* Wed Aug 05 09:20:39 2020



** Analysis setup **
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "complex_matlab_analysis.net"
.INC "complex_matlab_analysis.als"


.probe


.END
